`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.10.2022 15:06:45
// Design Name: 
// Module Name: cevrilebilir_and
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cevrilebilir_and(
    input A,B,
    output F
);
    cevrilebilir_kapi kullan(A,B,0,,F,);
endmodule
